`ifndef udp_uvm_include_pkg
`define udp_uvm_include_pkg

package udp_uvm_include_pkg;
	import uvm_pkg::*;
	`include "uvm_macros.svh"
	
	`include "udp_config.svh"
	`include "udp_transaction.svh"
	`include "udp_transaction.svh"
	`include "udp_sequences.svh"
	`include "udp_sequences.svh"
	`include "udp_virtual_sequences.svh"
	`include "udp_sequencer.svh"
	`include "udp_sequencer.svh"
	`include "udp_driver.svh"
	`include "udp_monitor.svh"
	`include "udp_driver.svh"
	`include "udp_monitor.svh"
	`include "udp_agent.svh"
	`include "udp_agent.svh"
	`include "udp_env.svh"
	`include "udp_tests.svh"
endpackage

import udp_uvm_include_pkg::*;

`endif