import global_typs_pkg::*;

module udp_vhdl_sv (
	udp_tx_if udp_tx_if_inst
	);

//Instance 
UDP_TX UDP_TX_inst (.*)


endmodule